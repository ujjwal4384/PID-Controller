`timescale 1ns / 1ps
//16 bit signed binary multiplier to give 16 bit output
module multiplier(A,B,ans);
input [15:0] A,B;
output [15:0]ans;
wire [31:0]M;
wire A0B0,A1B0,A2B0,A3B0,A4B0,A5B0,A6B0,A7B0,A8B0,A9B0,A10B0,A11B0,A12B0,A13B0,A14B0,A15B0;
wire A0B1,A1B1,A2B1,A3B1,A4B1,A5B1,A6B1,A7B1,A8B1,A9B1,A10B1,A11B1,A12B1,A13B1,A14B1,A15B1;
wire A0B2,A1B2,A2B2,A3B2,A4B2,A5B2,A6B2,A7B2,A8B2,A9B2,A10B2,A11B2,A12B2,A13B2,A14B2,A15B2;
wire A0B3,A1B3,A2B3,A3B3,A4B3,A5B3,A6B3,A7B3,A8B3,A9B3,A10B3,A11B3,A12B3,A13B3,A14B3,A15B3;
wire A0B4,A1B4,A2B4,A3B4,A4B4,A5B4,A6B4,A7B4,A8B4,A9B4,A10B4,A11B4,A12B4,A13B4,A14B4,A15B4;
wire A0B5,A1B5,A2B5,A3B5,A4B5,A5B5,A6B5,A7B5,A8B5,A9B5,A10B5,A11B5,A12B5,A13B5,A14B5,A15B5;
wire A0B6,A1B6,A2B6,A3B6,A4B6,A5B6,A6B6,A7B6,A8B6,A9B6,A10B6,A11B6,A12B6,A13B6,A14B6,A15B6;
wire A0B7,A1B7,A2B7,A3B7,A4B7,A5B7,A6B7,A7B7,A8B7,A9B7,A10B7,A11B7,A12B7,A13B7,A14B7,A15B7;
wire A0B8,A1B8,A2B8,A3B8,A4B8,A5B8,A6B8,A7B8,A8B8,A9B8,A10B8,A11B8,A12B8,A13B8,A14B8,A15B8;
wire A0B9,A1B9,A2B9,A3B9,A4B9,A5B9,A6B9,A7B9,A8B9,A9B9,A10B9,A11B9,A12B9,A13B9,A14B9,A15B9;
wire A0B10,A1B10,A2B10,A3B10,A4B10,A5B10,A6B10,A7B10,A8B10,A9B10,A10B10,A11B10,A12B10,A13B10,A14B10,A15B10;
wire A0B11,A1B11,A2B11,A3B11,A4B11,A5B11,A6B11,A7B11,A8B11,A9B11,A10B11,A11B11,A12B11,A13B11,A14B11,A15B11;
wire A0B12,A1B12,A2B12,A3B12,A4B12,A5B12,A6B12,A7B12,A8B12,A9B12,A10B12,A11B12,A12B12,A13B12,A14B12,A15B12;
wire A0B13,A1B13,A2B13,A3B13,A4B13,A5B13,A6B13,A7B13,A8B13,A9B13,A10B13,A11B13,A12B13,A13B13,A14B13,A15B13;
wire A0B14,A1B14,A2B14,A3B14,A4B14,A5B14,A6B14,A7B14,A8B14,A9B14,A10B14,A11B14,A12B14,A13B14,A14B14,A15B14;
wire A0B15,A1B15,A2B15,A3B15,A4B15,A5B15,A6B15,A7B15,A8B15,A9B15,A10B15,A11B15,A12B15,A13B15,A14B15,A15B15;
wire c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,temp;
wire [15:0] sum1,sum2,sum3,sum4,sum5,sum6,sum7,sum8,sum9,sum10,sum11,sum12,sum13,sum14,sum15;
wire [15:0] p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15;

and(A0B0,A[0],B[0]);
and(A1B0,A[1],B[0]);
and(A2B0,A[2],B[0]);
and(A3B0,A[3],B[0]);
and(A4B0,A[4],B[0]);
and(A5B0,A[5],B[0]);
and(A6B0,A[6],B[0]);
and(A7B0,A[7],B[0]);
and(A8B0,A[8],B[0]);
and(A9B0,A[9],B[0]);
and(A10B0,A[10],B[0]);
and(A11B0,A[11],B[0]);
and(A12B0,A[12],B[0]);
and(A13B0,A[13],B[0]);
and(A14B0,A[14],B[0]);
and(A15B0,A[15],B[0]);

and(A0B1,A[0],B[1]);
and(A1B1,A[1],B[1]);
and(A2B1,A[2],B[1]);
and(A3B1,A[3],B[1]);
and(A4B1,A[4],B[1]);
and(A5B1,A[5],B[1]);
and(A6B1,A[6],B[1]);
and(A7B1,A[7],B[1]);
and(A8B1,A[8],B[1]);
and(A9B1,A[9],B[1]);
and(A10B1,A[10],B[1]);
and(A11B1,A[11],B[1]);
and(A12B1,A[12],B[1]);
and(A13B1,A[13],B[1]);
and(A14B1,A[14],B[1]);
and(A15B1,A[15],B[1]);

and(A0B2,A[0],B[2]);
and(A1B2,A[1],B[2]);
and(A2B2,A[2],B[2]);
and(A3B2,A[3],B[2]);
and(A4B2,A[4],B[2]);
and(A5B2,A[5],B[2]);
and(A6B2,A[6],B[2]);
and(A7B2,A[7],B[2]);
and(A8B2,A[8],B[2]);
and(A9B2,A[9],B[2]);
and(A10B2,A[10],B[2]);
and(A11B2,A[11],B[2]);
and(A12B2,A[12],B[2]);
and(A13B2,A[13],B[2]);
and(A14B2,A[14],B[2]);
and(A15B2,A[15],B[2]);

and(A0B3,A[0],B[3]);
and(A1B3,A[1],B[3]);
and(A2B3,A[2],B[3]);
and(A3B3,A[3],B[3]);
and(A4B3,A[4],B[3]);
and(A5B3,A[5],B[3]);
and(A6B3,A[6],B[3]);
and(A7B3,A[7],B[3]);
and(A8B3,A[8],B[3]);
and(A9B3,A[9],B[3]);
and(A10B3,A[10],B[3]);
and(A11B3,A[11],B[3]);
and(A12B3,A[12],B[3]);
and(A13B3,A[13],B[3]);
and(A14B3,A[14],B[3]);
and(A15B3,A[15],B[3]);

and(A0B4,A[0],B[4]);
and(A1B4,A[1],B[4]);
and(A2B4,A[2],B[4]);
and(A3B4,A[3],B[4]);
and(A4B4,A[4],B[4]);
and(A5B4,A[5],B[4]);
and(A6B4,A[6],B[4]);
and(A7B4,A[7],B[4]);
and(A8B4,A[8],B[4]);
and(A9B4,A[9],B[4]);
and(A10B4,A[10],B[4]);
and(A11B4,A[11],B[4]);
and(A12B4,A[12],B[4]);
and(A13B4,A[13],B[4]);
and(A14B4,A[14],B[4]);
and(A15B4,A[15],B[4]);

and(A0B5,A[0],B[5]);
and(A1B5,A[1],B[5]);
and(A2B5,A[2],B[5]);
and(A3B5,A[3],B[5]);
and(A4B5,A[4],B[5]);
and(A5B5,A[5],B[5]);
and(A6B5,A[6],B[5]);
and(A7B5,A[7],B[5]);
and(A8B5,A[8],B[5]);
and(A9B5,A[9],B[5]);
and(A10B5,A[10],B[5]);
and(A11B5,A[11],B[5]);
and(A12B5,A[12],B[5]);
and(A13B5,A[13],B[5]);
and(A14B5,A[14],B[5]);
and(A15B5,A[15],B[5]);

and(A0B6,A[0],B[6]);
and(A1B6,A[1],B[6]);
and(A2B6,A[2],B[6]);
and(A3B6,A[3],B[6]);
and(A4B6,A[4],B[6]);
and(A5B6,A[5],B[6]);
and(A6B6,A[6],B[6]);
and(A7B6,A[7],B[6]);
and(A8B6,A[8],B[6]);
and(A9B6,A[9],B[6]);
and(A10B6,A[10],B[6]);
and(A11B6,A[11],B[6]);
and(A12B6,A[12],B[6]);
and(A13B6,A[13],B[6]);
and(A14B6,A[14],B[6]);
and(A15B6,A[15],B[6]);

and(A0B7,A[0],B[7]);
and(A1B7,A[1],B[7]);
and(A2B7,A[2],B[7]);
and(A3B7,A[3],B[7]);
and(A4B7,A[4],B[7]);
and(A5B7,A[5],B[7]);
and(A6B7,A[6],B[7]);
and(A7B7,A[7],B[7]);
and(A8B7,A[8],B[7]);
and(A9B7,A[9],B[7]);
and(A10B7,A[10],B[7]);
and(A11B7,A[11],B[7]);
and(A12B7,A[12],B[7]);
and(A13B7,A[13],B[7]);
and(A14B7,A[14],B[7]);
and(A15B7,A[15],B[7]);

and(A0B8,A[0],B[8]);
and(A1B8,A[1],B[8]);
and(A2B8,A[2],B[8]);
and(A3B8,A[3],B[8]);
and(A4B8,A[4],B[8]);
and(A5B8,A[5],B[8]);
and(A6B8,A[6],B[8]);
and(A7B8,A[7],B[8]);
and(A8B8,A[8],B[8]);
and(A9B8,A[9],B[8]);
and(A10B8,A[10],B[8]);
and(A11B8,A[11],B[8]);
and(A12B8,A[12],B[8]);
and(A13B8,A[13],B[8]);
and(A14B8,A[14],B[8]);
and(A15B8,A[15],B[8]);

and(A0B9,A[0],B[9]);
and(A1B9,A[1],B[9]);
and(A2B9,A[2],B[9]);
and(A3B9,A[3],B[9]);
and(A4B9,A[4],B[9]);
and(A5B9,A[5],B[9]);
and(A6B9,A[6],B[9]);
and(A7B9,A[7],B[9]);
and(A8B9,A[8],B[9]);
and(A9B9,A[9],B[9]);
and(A10B9,A[10],B[9]);
and(A11B9,A[11],B[9]);
and(A12B9,A[12],B[9]);
and(A13B9,A[13],B[9]);
and(A14B9,A[14],B[9]);
and(A15B9,A[15],B[9]);

and(A0B10,A[0],B[10]);
and(A1B10,A[1],B[10]);
and(A2B10,A[2],B[10]);
and(A3B10,A[3],B[10]);
and(A4B10,A[4],B[10]);
and(A5B10,A[5],B[10]);
and(A6B10,A[6],B[10]);
and(A7B10,A[7],B[10]);
and(A8B10,A[8],B[10]);
and(A9B10,A[9],B[10]);
and(A10B10,A[10],B[10]);
and(A11B10,A[11],B[10]);
and(A12B10,A[12],B[10]);
and(A13B10,A[13],B[10]);
and(A14B10,A[14],B[10]);
and(A15B10,A[15],B[10]);

and(A0B11,A[0],B[11]);
and(A1B11,A[1],B[11]);
and(A2B11,A[2],B[11]);
and(A3B11,A[3],B[11]);
and(A4B11,A[4],B[11]);
and(A5B11,A[5],B[11]);
and(A6B11,A[6],B[11]);
and(A7B11,A[7],B[11]);
and(A8B11,A[8],B[11]);
and(A9B11,A[9],B[11]);
and(A10B11,A[10],B[11]);
and(A11B11,A[11],B[11]);
and(A12B11,A[12],B[11]);
and(A13B11,A[13],B[11]);
and(A14B11,A[14],B[11]);
and(A15B11,A[15],B[11]);

and(A0B12,A[0],B[12]);
and(A1B12,A[1],B[12]);
and(A2B12,A[2],B[12]);
and(A3B12,A[3],B[12]);
and(A4B12,A[4],B[12]);
and(A5B12,A[5],B[12]);
and(A6B12,A[6],B[12]);
and(A7B12,A[7],B[12]);
and(A8B12,A[8],B[12]);
and(A9B12,A[9],B[12]);
and(A10B12,A[10],B[12]);
and(A11B12,A[11],B[12]);
and(A12B12,A[12],B[12]);
and(A13B12,A[13],B[12]);
and(A14B12,A[14],B[12]);
and(A15B12,A[15],B[12]);

and(A0B13,A[0],B[13]);
and(A1B13,A[1],B[13]);
and(A2B13,A[2],B[13]);
and(A3B13,A[3],B[13]);
and(A4B13,A[4],B[13]);
and(A5B13,A[5],B[13]);
and(A6B13,A[6],B[13]);
and(A7B13,A[7],B[13]);
and(A8B13,A[8],B[13]);
and(A9B13,A[9],B[13]);
and(A10B13,A[10],B[13]);
and(A11B13,A[11],B[13]);
and(A12B13,A[12],B[13]);
and(A13B13,A[13],B[13]);
and(A14B13,A[14],B[13]);
and(A15B13,A[15],B[13]);

and(A0B14,A[0],B[14]);
and(A1B14,A[1],B[14]);
and(A2B14,A[2],B[14]);
and(A3B14,A[3],B[14]);
and(A4B14,A[4],B[14]);
and(A5B14,A[5],B[14]);
and(A6B14,A[6],B[14]);
and(A7B14,A[7],B[14]);
and(A8B14,A[8],B[14]);
and(A9B14,A[9],B[14]);
and(A10B14,A[10],B[14]);
and(A11B14,A[11],B[14]);
and(A12B14,A[12],B[14]);
and(A13B14,A[13],B[14]);
and(A14B14,A[14],B[14]);
and(A15B14,A[15],B[14]);

and(A0B15,A[0],B[15]);
and(A1B15,A[1],B[15]);
and(A2B15,A[2],B[15]);
and(A3B15,A[3],B[15]);
and(A4B15,A[4],B[15]);
and(A5B15,A[5],B[15]);
and(A6B15,A[6],B[15]);
and(A7B15,A[7],B[15]);
and(A8B15,A[8],B[15]);
and(A9B15,A[9],B[15]);
and(A10B15,A[10],B[15]);
and(A11B15,A[11],B[15]);
and(A12B15,A[12],B[15]);
and(A13B15,A[13],B[15]);
and(A14B15,A[14],B[15]);
and(A15B15,A[15],B[15]);

buf(M[0],A0B0);
assign p0={1'b0,A15B0,A14B0,A13B0,A12B0,A11B0,A10B0,A9B0,A8B0,A7B0,A6B0,A5B0,A4B0,A3B0,A2B0,A1B0};
assign p1={A15B1,A14B1,A13B1,A12B1,A11B1,A10B1,A9B1,A8B1,A7B1,A6B1,A5B1,A4B1,A3B1,A2B1,A1B1,A0B1};
assign p2={A15B2,A14B2,A13B2,A12B2,A11B2,A10B2,A9B2,A8B2,A7B2,A6B2,A5B2,A4B2,A3B2,A2B2,A1B2,A0B2};
assign p3={A15B3,A14B3,A13B3,A12B3,A11B3,A10B3,A9B3,A8B3,A7B3,A6B3,A5B3,A4B3,A3B3,A2B3,A1B3,A0B3};
assign p4={A15B4,A14B4,A13B4,A12B4,A11B4,A10B4,A9B4,A8B4,A7B4,A6B4,A5B4,A4B4,A3B4,A2B4,A1B4,A0B4};
assign p5={A15B5,A14B5,A13B5,A12B5,A11B5,A10B5,A9B5,A8B5,A7B5,A6B5,A5B5,A4B5,A3B5,A2B5,A1B5,A0B5};
assign p6={A15B6,A14B6,A13B6,A12B6,A11B6,A10B6,A9B6,A8B6,A7B6,A6B6,A5B6,A4B6,A3B6,A2B6,A1B6,A0B6};
assign p7={A15B7,A14B7,A13B7,A12B7,A11B7,A10B7,A9B7,A8B7,A7B7,A6B7,A5B7,A4B7,A3B7,A2B7,A1B7,A0B7};
assign p8={A15B8,A14B8,A13B8,A12B8,A11B8,A10B8,A9B8,A8B8,A7B8,A6B8,A5B8,A4B8,A3B8,A2B8,A1B8,A0B8};
assign p9={A15B9,A14B9,A13B9,A12B9,A11B9,A10B9,A9B9,A8B9,A7B9,A6B9,A5B9,A4B9,A3B9,A2B9,A1B9,A0B9};
assign p10={A15B10,A14B10,A13B10,A12B10,A11B10,A10B10,A9B10,A8B10,A7B10,A6B10,A5B10,A4B10,A3B10,A2B10,A1B10,A0B10};
assign p11={A15B11,A14B11,A13B11,A12B11,A11B11,A10B11,A9B11,A8B11,A7B11,A6B11,A5B11,A4B11,A3B11,A2B11,A1B11,A0B11};
assign p12={A15B12,A14B12,A13B12,A12B12,A11B12,A10B12,A9B12,A8B12,A7B12,A6B12,A5B12,A4B12,A3B12,A2B12,A1B12,A0B12};
assign p13={A15B13,A14B13,A13B13,A12B13,A11B13,A10B13,A9B13,A8B13,A7B13,A6B13,A5B13,A4B13,A3B13,A2B13,A1B13,A0B13};
assign p14={A15B14,A14B14,A13B14,A12B14,A11B14,A10B14,A9B14,A8B14,A7B14,A6B14,A5B14,A4B14,A3B14,A2B14,A1B14,A0B14};
assign p15={A15B15,A14B15,A13B15,A12B15,A11B15,A10B15,A9B15,A8B15,A7B15,A6B15,A5B15,A4B15,A3B15,A2B15,A1B15,A0B15};

_16BitAdder A0(p0,p1,1'b0,sum1,c1);
buf(M[1],sum1[0]);
_16BitAdder A1({c1,sum1[15:1]},p2,1'b0,sum2,c2);
buf(M[2],sum2[0]);
_16BitAdder A2({c2,sum2[15:1]},p3,1'b0,sum3,c3);
buf(M[3],sum3[0]);
_16BitAdder A3({c3,sum3[15:1]},p4,1'b0,sum4,c4);
buf(M[4],sum4[0]);
_16BitAdder A4({c4,sum4[15:1]},p5,1'b0,sum5,c5);
buf(M[5],sum5[0]);
_16BitAdder A5({c5,sum5[15:1]},p6,1'b0,sum6,c6);
buf(M[6],sum6[0]);
_16BitAdder A6({c6,sum6[15:1]},p7,1'b0,sum7,c7);
buf(M[7],sum7[0]);
_16BitAdder A7({c7,sum7[15:1]},p8,1'b0,sum8,c8);
buf(M[8],sum8[0]);
_16BitAdder A8({c8,sum8[15:1]},p9,1'b0,sum9,c9);
buf(M[9],sum9[0]);
_16BitAdder A9({c9,sum9[15:1]},p10,1'b0,sum10,c10);
buf(M[10],sum10[0]);
_16BitAdder A10({c10,sum10[15:1]},p11,1'b0,sum11,c11);
buf(M[11],sum11[0]);
_16BitAdder A11({c11,sum11[15:1]},p12,1'b0,sum12,c12);
buf(M[12],sum12[0]);
_16BitAdder A12({c12,sum12[15:1]},p13,1'b0,sum13,c13);
buf(M[13],sum13[0]);
_16BitAdder A13({c13,sum13[15:1]},p14,1'b0,sum14,c14);
buf(M[14],sum14[0]);
_16BitAdder A14({c14,sum14[15:1]},p15,1'b0,sum15,c15);
assign ans={sum15[0],M[14:0]};
endmodule